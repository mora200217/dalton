// Sumador.v

module sum(
               input a,
               input b,
               output c
               );


   assign c = a & b;

endmodule // prueba
